`ifndef LSU_VH
`define LSU_VH

`define LSUOP_WIDTH 3
`define LSUOP_B    `LSUOP_WIDTH'd00
`define LSUOP_H    `LSUOP_WIDTH'd01
`define LSUOP_W    `LSUOP_WIDTH'd02
`define LSUOP_BU   `LSUOP_WIDTH'd03
`define LSUOP_HU   `LSUOP_WIDTH'd04
`define LSUOP_X    `LSUOP_WIDTH'dX

`endif
